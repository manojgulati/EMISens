* C:\Users\Omkar\Dropbox\EMI_Sense_Design_project\PSpice_simulations\ver1.6\Differential_filter(680Vpp)_test_18_march.sch

* Schematics Version 9.1 - Web Update 1
* Wed Mar 26 14:57:49 2014



** Analysis setup **
.ac LIN 10001 1 10000.00K
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Differential_filter(680Vpp)_test_18_march.net"
.INC "Differential_filter(680Vpp)_test_18_march.als"


.probe


.END
