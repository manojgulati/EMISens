* C:\Users\manojg\Dropbox\EMI_Sense_Design_project\PSpice_simulations\ver1.5\Schematic2.sch

* Schematics Version 9.1 - Web Update 1
* Sat Mar 01 17:08:52 2014



** Analysis setup **
.ac LIN 101 10 500.00K
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic2.net"
.INC "Schematic2.als"


.probe


.END
