* C:\Users\manojg\Dropbox\EMI_Sense_Design_project\PSpice_simulations\ver1.2\Filter_ver1.2.sch

* Schematics Version 9.1 - Web Update 1
* Wed Jan 29 12:35:15 2014



** Analysis setup **
.ac LIN 101 10 500.00K
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Filter_ver1.2.net"
.INC "Filter_ver1.2.als"


.probe


.END
