* C:\Users\manojg\Dropbox\EMI_Sense_Design_project\PSpice_simulations\ver1.6\Schematic1.sch

* Schematics Version 9.1 - Web Update 1
* Sun Mar 02 15:18:22 2014



** Analysis setup **
.ac LIN 101 10 100.00K
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic1.net"
.INC "Schematic1.als"


.probe


.END
