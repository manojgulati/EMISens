* C:\Users\manojg\Dropbox\EMI_Sense_Design_project\PSpice_simulations\ver1.3\Schematic3.sch

* Schematics Version 9.1 - Web Update 1
* Tue Feb 18 21:55:34 2014



** Analysis setup **
.ac LIN 101 1K 500.00K
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic3.net"
.INC "Schematic3.als"


.probe


.END
