* C:\Users\manojg\Dropbox\EMI_Sense_Design_project\PSpice_simulations\ver1.4\Schematic1.sch

* Schematics Version 9.1 - Web Update 1
* Tue Feb 25 22:55:26 2014



** Analysis setup **
.ac LIN 101 10 1.00K
.tran 10ms 100s
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic1.net"
.INC "Schematic1.als"


.probe


.END
