* C:\Users\manojg\Dropbox\EMI_Sense_Design_project\PSpice_simulations\ver1.5\Schematic5.sch

* Schematics Version 9.1 - Web Update 1
* Sat Mar 01 11:39:05 2014



** Analysis setup **
.ac LIN 101 10 100.00K
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic5.net"
.INC "Schematic5.als"


.probe


.END
