* C:\Users\manojg\Dropbox\EMI_Sense_Design_project\PSpice_simulations\ver1.3\Schematic6.sch

* Schematics Version 9.1 - Web Update 1
* Wed Feb 19 22:30:01 2014



** Analysis setup **
.ac LIN 100 100 1000.00K
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic6.net"
.INC "Schematic6.als"


.probe


.END
