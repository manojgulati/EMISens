* C:\Users\Omkar\Dropbox\EMI_Sense_Design_project\PSpice_simulations\ver1.2\Filter_ver1.3.sch

* Schematics Version 9.1 - Web Update 1
* Mon Feb 03 23:31:59 2014



** Analysis setup **
.ac LIN 101 10 500.00K
.tran 0ns 1000ns
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Filter_ver1.3.net"
.INC "Filter_ver1.3.als"


.probe


.END
