* C:\Users\Omkar\Dropbox\EMI_Sense_Design_project\PSpice_simulations\ver1.4\FLT_6.sch

* Schematics Version 9.1 - Web Update 1
* Sat Feb 22 01:03:42 2014



** Analysis setup **
.ac LIN 101 10 350.00K
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "FLT_6.net"
.INC "FLT_6.als"


.probe


.END
