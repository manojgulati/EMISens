* C:\Users\manojg\Dropbox\EMI_Sense_Design_project\PSpice_simulations\ver1.3\Schematic4.sch

* Schematics Version 9.1 - Web Update 1
* Tue Feb 18 23:19:41 2014



** Analysis setup **
.ac LIN 101 1K 500.00K
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic4.net"
.INC "Schematic4.als"


.probe


.END
