* C:\Users\manojg\Dropbox\EMI_Sense_Design_project\PSpice_simulations\ver1.6\Differential_filter(680Vpp).sch

* Schematics Version 9.1 - Web Update 1
* Mon Mar 03 21:50:52 2014



** Analysis setup **
.ac LIN 101 10 400.00K
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Differential_filter(680Vpp).net"
.INC "Differential_filter(680Vpp).als"


.probe


.END
