* C:\Users\manojg\Dropbox\EMI_Sense_Design_project\PSpice_simulations\Filter_ver1.1.sch

* Schematics Version 9.1 - Web Update 1
* Wed Jan 29 12:04:50 2014



** Analysis setup **
.ac LIN 101 10 250.00K
.tran 0ns 1000ns
.OP 
.STMLIB "Filter_ver1.1.stl"


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Filter_ver1.1.net"
.INC "Filter_ver1.1.als"


.probe


.END
