* C:\Users\Omkar\Dropbox\EMI_Sense_Design_project\PSpice_simulations\ver1.2\Filter_ver1.4.sch

* Schematics Version 9.1 - Web Update 1
* Mon Feb 03 23:39:49 2014



** Analysis setup **
.ac LIN 101 10 500.00K
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Filter_ver1.4.net"
.INC "Filter_ver1.4.als"


.probe


.END
