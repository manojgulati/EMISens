* C:\Users\Omkar\Dropbox\EMI_Sense_Design_project\PSpice_simulations\ver1.6\Differential_filter(680Vpp)_Power_test.sch

* Schematics Version 9.1 - Web Update 1
* Fri Mar 07 11:53:31 2014



** Analysis setup **
.tran/OP 0ns 1000ns
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Differential_filter(680Vpp)_Power_test.net"
.INC "Differential_filter(680Vpp)_Power_test.als"


.probe


.END
