* C:\Users\manojg\Dropbox\EMI_Sense_Design_project\PSpice_simulations\ver1.6\Differential_filter(680Vpp)_test.sch

* Schematics Version 9.1 - Web Update 1
* Mon Mar 03 23:37:45 2014



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Differential_filter(680Vpp)_test.net"
.INC "Differential_filter(680Vpp)_test.als"


.probe


.END
