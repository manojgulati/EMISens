* C:\Users\Omkar\Dropbox\EMI_Sense_Design_project\PSpice_simulations\ver1.6\Differential_filter(680Vpp)_test_2.sch

* Schematics Version 9.1 - Web Update 1
* Tue Mar 04 20:15:58 2014



** Analysis setup **
.ac LIN 101 10 2000.00K
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Differential_filter(680Vpp)_test_2.net"
.INC "Differential_filter(680Vpp)_test_2.als"


.probe


.END
