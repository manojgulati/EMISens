* C:\Users\manojg\Dropbox\EMI_Sense_Design_project\PSpice_simulations\ver1.3\Schematic1.sch

* Schematics Version 9.1 - Web Update 1
* Tue Feb 18 20:59:33 2014



** Analysis setup **
.ac LIN 101 1K 350.00K
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic1.net"
.INC "Schematic1.als"


.probe


.END
